`timescale 1ns/100ps

module mult255 (
   input iclk,
   input irst_n,

   input      [7:0]  x,
   output reg [15:0] q
);

   `ifdef COCOTB_SIM
    initial begin
      $dumpfile("mult255_wave.vcd");
      $dumpvars(0, mult255);
      #1;
    end
  `endif

   always @(posedge iclk) begin
      if (!irst_n)
         q <= 16'h0000;
      else begin
         case (x)
            8'h00 : q <= 16'h0000;
            8'h01 : q <= 16'h00ff;
            8'h02 : q <= 16'h01fe;
            8'h03 : q <= 16'h02fd;
            8'h04 : q <= 16'h03fc;
            8'h05 : q <= 16'h04fb;
            8'h06 : q <= 16'h05fa;
            8'h07 : q <= 16'h06f9;
            8'h08 : q <= 16'h07f8;
            8'h09 : q <= 16'h08f7;
            8'h0A : q <= 16'h09f6;
            8'h0B : q <= 16'h0af5;
            8'h0C : q <= 16'h0bf4;
            8'h0D : q <= 16'h0cf3;
            8'h0E : q <= 16'h0df2;
            8'h0F : q <= 16'h0ef1;
            8'h10 : q <= 16'h0ff0;
            8'h11 : q <= 16'h10ef;
            8'h12 : q <= 16'h11ee;
            8'h13 : q <= 16'h12ed;
            8'h14 : q <= 16'h13ec;
            8'h15 : q <= 16'h14eb;
            8'h16 : q <= 16'h15ea;
            8'h17 : q <= 16'h16e9;
            8'h18 : q <= 16'h17e8;
            8'h19 : q <= 16'h18e7;
            8'h1A : q <= 16'h19e6;
            8'h1B : q <= 16'h1ae5;
            8'h1C : q <= 16'h1be4;
            8'h1D : q <= 16'h1ce3;
            8'h1E : q <= 16'h1de2;
            8'h1F : q <= 16'h1ee1;
            8'h20 : q <= 16'h1fe0;
            8'h21 : q <= 16'h20df;
            8'h22 : q <= 16'h21de;
            8'h23 : q <= 16'h22dd;
            8'h24 : q <= 16'h23dc;
            8'h25 : q <= 16'h24db;
            8'h26 : q <= 16'h25da;
            8'h27 : q <= 16'h26d9;
            8'h28 : q <= 16'h27d8;
            8'h29 : q <= 16'h28d7;
            8'h2A : q <= 16'h29d6;
            8'h2B : q <= 16'h2ad5;
            8'h2C : q <= 16'h2bd4;
            8'h2D : q <= 16'h2cd3;
            8'h2E : q <= 16'h2dd2;
            8'h2F : q <= 16'h2ed1;
            8'h30 : q <= 16'h2fd0;
            8'h31 : q <= 16'h30cf;
            8'h32 : q <= 16'h31ce;
            8'h33 : q <= 16'h32cd;
            8'h34 : q <= 16'h33cc;
            8'h35 : q <= 16'h34cb;
            8'h36 : q <= 16'h35ca;
            8'h37 : q <= 16'h36c9;
            8'h38 : q <= 16'h37c8;
            8'h39 : q <= 16'h38c7;
            8'h3A : q <= 16'h39c6;
            8'h3B : q <= 16'h3ac5;
            8'h3C : q <= 16'h3bc4;
            8'h3D : q <= 16'h3cc3;
            8'h3E : q <= 16'h3dc2;
            8'h3F : q <= 16'h3ec1;
            8'h40 : q <= 16'h3fc0;
            8'h41 : q <= 16'h40bf;
            8'h42 : q <= 16'h41be;
            8'h43 : q <= 16'h42bd;
            8'h44 : q <= 16'h43bc;
            8'h45 : q <= 16'h44bb;
            8'h46 : q <= 16'h45ba;
            8'h47 : q <= 16'h46b9;
            8'h48 : q <= 16'h47b8;
            8'h49 : q <= 16'h48b7;
            8'h4A : q <= 16'h49b6;
            8'h4B : q <= 16'h4ab5;
            8'h4C : q <= 16'h4bb4;
            8'h4D : q <= 16'h4cb3;
            8'h4E : q <= 16'h4db2;
            8'h4F : q <= 16'h4eb1;
            8'h50 : q <= 16'h4fb0;
            8'h51 : q <= 16'h50af;
            8'h52 : q <= 16'h51ae;
            8'h53 : q <= 16'h52ad;
            8'h54 : q <= 16'h53ac;
            8'h55 : q <= 16'h54ab;
            8'h56 : q <= 16'h55aa;
            8'h57 : q <= 16'h56a9;
            8'h58 : q <= 16'h57a8;
            8'h59 : q <= 16'h58a7;
            8'h5A : q <= 16'h59a6;
            8'h5B : q <= 16'h5aa5;
            8'h5C : q <= 16'h5ba4;
            8'h5D : q <= 16'h5ca3;
            8'h5E : q <= 16'h5da2;
            8'h5F : q <= 16'h5ea1;
            8'h60 : q <= 16'h5fa0;
            8'h61 : q <= 16'h609f;
            8'h62 : q <= 16'h619e;
            8'h63 : q <= 16'h629d;
            8'h64 : q <= 16'h639c;
            8'h65 : q <= 16'h649b;
            8'h66 : q <= 16'h659a;
            8'h67 : q <= 16'h6699;
            8'h68 : q <= 16'h6798;
            8'h69 : q <= 16'h6897;
            8'h6A : q <= 16'h6996;
            8'h6B : q <= 16'h6a95;
            8'h6C : q <= 16'h6b94;
            8'h6D : q <= 16'h6c93;
            8'h6E : q <= 16'h6d92;
            8'h6F : q <= 16'h6e91;
            8'h70 : q <= 16'h6f90;
            8'h71 : q <= 16'h708f;
            8'h72 : q <= 16'h718e;
            8'h73 : q <= 16'h728d;
            8'h74 : q <= 16'h738c;
            8'h75 : q <= 16'h748b;
            8'h76 : q <= 16'h758a;
            8'h77 : q <= 16'h7689;
            8'h78 : q <= 16'h7788;
            8'h79 : q <= 16'h7887;
            8'h7A : q <= 16'h7986;
            8'h7B : q <= 16'h7a85;
            8'h7C : q <= 16'h7b84;
            8'h7D : q <= 16'h7c83;
            8'h7E : q <= 16'h7d82;
            8'h7F : q <= 16'h7e81;
            8'h80 : q <= 16'h7f80;
            8'h81 : q <= 16'h807f;
            8'h82 : q <= 16'h817e;
            8'h83 : q <= 16'h827d;
            8'h84 : q <= 16'h837c;
            8'h85 : q <= 16'h847b;
            8'h86 : q <= 16'h857a;
            8'h87 : q <= 16'h8679;
            8'h88 : q <= 16'h8778;
            8'h89 : q <= 16'h8877;
            8'h8A : q <= 16'h8976;
            8'h8B : q <= 16'h8a75;
            8'h8C : q <= 16'h8b74;
            8'h8D : q <= 16'h8c73;
            8'h8E : q <= 16'h8d72;
            8'h8F : q <= 16'h8e71;
            8'h90 : q <= 16'h8f70;
            8'h91 : q <= 16'h906f;
            8'h92 : q <= 16'h916e;
            8'h93 : q <= 16'h926d;
            8'h94 : q <= 16'h936c;
            8'h95 : q <= 16'h946b;
            8'h96 : q <= 16'h956a;
            8'h97 : q <= 16'h9669;
            8'h98 : q <= 16'h9768;
            8'h99 : q <= 16'h9867;
            8'h9A : q <= 16'h9966;
            8'h9B : q <= 16'h9a65;
            8'h9C : q <= 16'h9b64;
            8'h9D : q <= 16'h9c63;
            8'h9E : q <= 16'h9d62;
            8'h9F : q <= 16'h9e61;
            8'hA0 : q <= 16'h9f60;
            8'hA1 : q <= 16'ha05f;
            8'hA2 : q <= 16'ha15e;
            8'hA3 : q <= 16'ha25d;
            8'hA4 : q <= 16'ha35c;
            8'hA5 : q <= 16'ha45b;
            8'hA6 : q <= 16'ha55a;
            8'hA7 : q <= 16'ha659;
            8'hA8 : q <= 16'ha758;
            8'hA9 : q <= 16'ha857;
            8'hAA : q <= 16'ha956;
            8'hAB : q <= 16'haa55;
            8'hAC : q <= 16'hab54;
            8'hAD : q <= 16'hac53;
            8'hAE : q <= 16'had52;
            8'hAF : q <= 16'hae51;
            8'hB0 : q <= 16'haf50;
            8'hB1 : q <= 16'hb04f;
            8'hB2 : q <= 16'hb14e;
            8'hB3 : q <= 16'hb24d;
            8'hB4 : q <= 16'hb34c;
            8'hB5 : q <= 16'hb44b;
            8'hB6 : q <= 16'hb54a;
            8'hB7 : q <= 16'hb649;
            8'hB8 : q <= 16'hb748;
            8'hB9 : q <= 16'hb847;
            8'hBA : q <= 16'hb946;
            8'hBB : q <= 16'hba45;
            8'hBC : q <= 16'hbb44;
            8'hBD : q <= 16'hbc43;
            8'hBE : q <= 16'hbd42;
            8'hBF : q <= 16'hbe41;
            8'hC0 : q <= 16'hbf40;
            8'hC1 : q <= 16'hc03f;
            8'hC2 : q <= 16'hc13e;
            8'hC3 : q <= 16'hc23d;
            8'hC4 : q <= 16'hc33c;
            8'hC5 : q <= 16'hc43b;
            8'hC6 : q <= 16'hc53a;
            8'hC7 : q <= 16'hc639;
            8'hC8 : q <= 16'hc738;
            8'hC9 : q <= 16'hc837;
            8'hCA : q <= 16'hc936;
            8'hCB : q <= 16'hca35;
            8'hCC : q <= 16'hcb34;
            8'hCD : q <= 16'hcc33;
            8'hCE : q <= 16'hcd32;
            8'hCF : q <= 16'hce31;
            8'hD0 : q <= 16'hcf30;
            8'hD1 : q <= 16'hd02f;
            8'hD2 : q <= 16'hd12e;
            8'hD3 : q <= 16'hd22d;
            8'hD4 : q <= 16'hd32c;
            8'hD5 : q <= 16'hd42b;
            8'hD6 : q <= 16'hd52a;
            8'hD7 : q <= 16'hd629;
            8'hD8 : q <= 16'hd728;
            8'hD9 : q <= 16'hd827;
            8'hDA : q <= 16'hd926;
            8'hDB : q <= 16'hda25;
            8'hDC : q <= 16'hdb24;
            8'hDD : q <= 16'hdc23;
            8'hDE : q <= 16'hdd22;
            8'hDF : q <= 16'hde21;
            8'hE0 : q <= 16'hdf20;
            8'hE1 : q <= 16'he01f;
            8'hE2 : q <= 16'he11e;
            8'hE3 : q <= 16'he21d;
            8'hE4 : q <= 16'he31c;
            8'hE5 : q <= 16'he41b;
            8'hE6 : q <= 16'he51a;
            8'hE7 : q <= 16'he619;
            8'hE8 : q <= 16'he718;
            8'hE9 : q <= 16'he817;
            8'hEA : q <= 16'he916;
            8'hEB : q <= 16'hea15;
            8'hEC : q <= 16'heb14;
            8'hED : q <= 16'hec13;
            8'hEE : q <= 16'hed12;
            8'hEF : q <= 16'hee11;
            8'hF0 : q <= 16'hef10;
            8'hF1 : q <= 16'hf00f;
            8'hF2 : q <= 16'hf10e;
            8'hF3 : q <= 16'hf20d;
            8'hF4 : q <= 16'hf30c;
            8'hF5 : q <= 16'hf40b;
            8'hF6 : q <= 16'hf50a;
            8'hF7 : q <= 16'hf609;
            8'hF8 : q <= 16'hf708;
            8'hF9 : q <= 16'hf807;
            8'hFA : q <= 16'hf906;
            8'hFB : q <= 16'hfa05;
            8'hFC : q <= 16'hfb04;
            8'hFD : q <= 16'hfc03;
            8'hFE : q <= 16'hfd02;
            8'hFF : q <= 16'hfe01;
            
            default : q <= 16'h0000;
         endcase
      end
   end

endmodule
